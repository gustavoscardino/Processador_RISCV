module rom64x32 (
    input [5:0] endereco,
    input clk,
    output [31:0] saida
);

     reg [32:0] rom [63:0];
     
    initial begin
        rom[0]   =   {12'd1 , 5'd0 , 3'b010 , 5'd1 , 7'b0000011}; // lw x1,x0(1)
        rom[4]   =   {12'd2 , 5'd0 , 3'b010 , 5'd2 , 7'b0000011}; //lw x2,x0(2)
        rom[8]   =   {12'd3 , 5'd0 , 3'b010 , 5'd3 , 7'b0000011}; //lw x3,x0(3)
        rom[12]  =   {}


        end


   assign saida = rom[endereco];

endmodule


//Instrucoes antigas
        //             rom[0]=  {12'd1 , 5'd0 , 3'b010 , 5'd1 , 7'b0000011}; // lw x1,x0(1)
        //             rom[4]=  {12'd2 , 5'd0 , 3'b010 , 5'd2 , 7'b0000011}; //lw x2,x0(2)
        //             rom[8]=  {12'd3 , 5'd0 , 3'b010 , 5'd3 , 7'b0000011}; //lw x3,x0(3)
        // /*while*/   rom[12]= {7'b0000001, 5'd2, 5'd1, 3'b000, 5'b00000, 7'b1100011}; //beq x1,x2,fim(+32)
        //             rom[16]= {7'b0100000, 5'd2, 5'd1, 3'b000, 5'd5, 7'b0110011}; //sub x5,x1,x2
        //             rom[20]= {7'b0000000, 5'd3, 5'd5, 3'b111, 5'd6, 7'b0110011}; //and x6, x5, x3
        //             rom[24]= {7'b0000000, 5'd3, 5'd6, 3'b000, 5'b01100, 7'b1100011}; //beq x6, x3, m(+12)
        //             rom[28]= {7'b0100000, 5'd2, 5'd1, 3'b000, 5'b1, 7'b0110011}; //sub x1,x1,x2 
        //             rom[32]= {7'b1111111, 5'd0, 5'd0, 3'b000, 5'b01101, 7'b1100011}; //beq x0,x0,while (-20)
        // /*m*/       rom[36]= {7'b0100000, 5'd1, 5'd2, 3'b000, 5'd2, 7'b0110011}; //sub x2,x2,x1
        //             rom[40]= {7'b0100000, 5'd0, 5'd0, 3'b000, 5'd2, 7'b0110011}; //beq x0,x0,while (-28)
        // /*fim*/     rom[44]= {7'b0000000, 5'd1, 5'd0, 3'b010, 5'b01010, 7'b0000011}; //sw x1,x0(10)